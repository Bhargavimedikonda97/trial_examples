module comb(comb_in, comb_out);
  input comb_in;
  output logic comb_out;
  assign comb_out = comb_in;
  endmodule
